`ifndef vertexinput_DEFINES
`define vertexinput_DEFINES

`define ADDR_W 32
`define DATA_W 32
`define BYTE 8
`define DATA_W_BYTES `DATA_W/`BYTE
`define NUMBER_REGISTERS 2

`endif
